module NOT(Y,A);
	input A;
	output Y;
	nand(Y,A,A);
endmodule
