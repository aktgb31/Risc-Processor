module D_FLIP_FLOP_FE_SR(Q,Q_,D,CLK,R);
    input D,CLK,R;
    output Q,Q_;
    wire r,d;
    nand(r,R,R);
    AND and_1(d,D,r);
    D_FLIP_FLOP_RE d1(Q,Q_,d,CLK);

endmodule

module D_FLIP_FLOP_FE(Q,Q_,D,CLK);
    input D,CLK;
    output Q,Q_;
    wire c,q;
    nand(c,CLK,CLK);
    D_LATCH d1(q,,D,CLK);
    D_LATCH d2(Q,Q_,q,c);

endmodule

module D_LATCH(Q,Q_,D,CLK);
    input D,CLK;
    output Q,Q_;
    wire a,b;
    nand(a,D,CLK);
    nand(b,a,CLK);
    nand(Q,Q_,a);
    nand(Q_,Q,b);
endmodule

module AND(Y,A,B);
	input A,B;
	output Y;
	wire x;	
	nand(x,A,B);
	nand(Y,x,x);
endmodule


